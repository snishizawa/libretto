* Library name: sg13g2_stdcell
* Cell name: sg13g2_o21ai_1
* View name: schematic
* Inherited view list: spectre cmos_sch cmos.sch schematic veriloga ahdl
* pspice dspf
.subckt sg13g2_o21ai_1 A1 A2 B1 VDD VSS Y
XP2 net14 A1 VDD VDD sg13_lv_pmos w=1.12u l=150.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XP1 Y A2 net14 VDD sg13_lv_pmos w=1.12u l=150.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XP0 Y B1 VDD VDD sg13_lv_pmos w=1.12u l=150.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XN2 net1 A2 VSS VSS sg13_lv_nmos w=740.00n l=150.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XN3 net1 A1 VSS VSS sg13_lv_nmos w=740.00n l=150.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XN0 Y B1 net1 VSS sg13_lv_nmos w=740.00n l=150.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
.ends
* End of subcircuit definition.
