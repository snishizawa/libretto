.subckt AO22_1X A1 A2 B1 B2 Y VDD VSS VNW VPW
MP1 VDD A1 w1  VNW p m=1 L=350n W=1800n
MP2 VDD A2 w1  VNW p m=1 L=350n W=1800n
MP3 w1  B1 YB  VNW p m=1 L=350n W=1800n
MP4 w1  B2 YB  VNW p m=1 L=350n W=1800n
MN1 VSS A1 w2  VPW n m=1 L=350n W=1200n
MN2 w2  A2 YB  VPW n m=1 L=350n W=1200n
MN3 VSS B1 w3  VPW n m=1 L=350n W=1200n
MN4 w3  B2 YB  VPW n m=1 L=350n W=1200n
MP5 VDD YB Y VNW p m=1 L=350n W=1800n
MN5 VSS YB Y VPW n m=1 L=350n W=1200n
.ends
