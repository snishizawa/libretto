* Library name: sg13g2_stdcell
* Cell name: sg13g2_nor2_2
* View name: schematic
* Inherited view list: spectre cmos_sch cmos.sch schematic veriloga ahdl
* pspice dspf
.subckt sg13g2_nor2_2 A B VDD VSS Y
XX0 Y A VSS VSS sg13_lv_nmos w=1.48u l=130.00n ng=2 ad=0 as=0 pd=0 ps=0 m=1
XX3 Y B VSS VSS sg13_lv_nmos w=1.48u l=130.00n ng=2 ad=0 as=0 pd=0 ps=0 m=1
XX1 net1 A VDD VDD sg13_lv_pmos w=2.24u l=130.00n ng=2 ad=0 as=0 pd=0 ps=0 m=1
XX2 Y B net1 VDD sg13_lv_pmos w=2.24u l=130.00n ng=2 ad=0 as=0 pd=0 ps=0 m=1
.ends
* End of subcircuit definition.
