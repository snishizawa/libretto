.subckt OR4_1X A B C D Y VDD VSS VNW VPW
MP1 VDD A W1 VNW p m=1 L=350n W=1800n
MP2 W1  B W2 VNW p m=1 L=350n W=1800n
MP3 W2  C W3 VNW p m=1 L=350n W=1800n
MP4 W3  D YB VNW p m=1 L=350n W=1800n
MN1 VSS A YB VPW n m=1 L=350n W=1200n
MN2 VSS B YB VPW n m=1 L=350n W=1200n
MN3 VSS C YB VPW n m=1 L=350n W=1200n
MN4 VSS D YB VPW n m=1 L=350n W=1200n
MP5 VDD YB Y VNW p m=1 L=350n W=1800n
MN5 VSS YB Y VPW n m=1 L=350n W=1200n
.ends
