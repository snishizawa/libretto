* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_isobufsrc_8 A SLEEP VGND VNB VPB VPWR X
X0 a_321_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_123_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 X a_123_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A a_123_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_123_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_123_297# a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_321_297# a_123_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 X a_123_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_321_297# a_123_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_321_297# a_123_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_321_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_321_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR a_123_297# a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 X a_123_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 X SLEEP a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_123_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 X SLEEP a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VGND a_123_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VGND A a_123_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VGND a_123_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VGND a_123_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VPWR a_123_297# a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VPWR a_123_297# a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 a_123_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 X SLEEP a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 X SLEEP a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 a_321_297# a_123_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 a_321_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends
