.subckt OR2_1X A B Y VDD VSS VNW VPW
MP1 VDD A W1 VNW p m=1    L=350n W=1800n
MP2 W1  B YB VNW p m=1    L=350n W=1800n
MN1 VSS A YB VPW n m=1    L=350n W=1200n
MN2 VSS B YB VPW n m=1    L=350n W=1200n
MP3 VDD YB Y VNW p m=1 L=350n W=1800n
MN3 VSS YB Y VPW n m=1 L=350n W=1200n
.ends
