* Library name: sg13g2_stdcell
* Cell name: sg13g2_nor3_1
* View name: schematic
* Inherited view list: spectre cmos_sch cmos.sch schematic veriloga ahdl
* pspice dspf
.subckt sg13g2_nor3_1 A B C VDD VSS Y
XX3 net1 C Y VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX0 net2 B net1 VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX2 VDD A net2 VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX4 Y A VSS VSS sg13_lv_nmos w=770.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX1 Y B VSS VSS sg13_lv_nmos w=770.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX5 Y C VSS VSS sg13_lv_nmos w=770.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
.ends
* End of subcircuit definition.
