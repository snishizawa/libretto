* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_471_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_1241_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_297# B1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_471_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_27_297# B1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND A2 a_1241_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_471_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_453_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_471_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_471_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 Y A1 a_1241_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND A2 a_1241_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VGND B2 a_453_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_471_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VGND B2 a_453_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_453_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR A1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 VPWR A1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_453_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_1241_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 a_1241_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_27_297# B2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 VPWR A2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_471_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 a_1241_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 a_471_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 VPWR A2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 Y B1 a_453_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 a_27_297# B2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X37 Y B1 a_453_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 Y A1 a_1241_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 a_453_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
