.subckt XNOR2_1X A B Y VDD VSS VNW VPW
* AINV
MP1 VDD A AB VNW p m=1 L=350n W=1800n
MN1 VSS A AB VPW n m=1 L=350n W=1200n

* BINV
MP2 VDD B BB VNW p m=1 L=350n W=1800n
MN2 VSS B BB VPW n m=1 L=350n W=1200n

* TGB
MP3 B A  TG VNW p m=1 L=350n W=1800n
MN3 B AB TG VPW n m=1 L=350n W=1200n

* TGBB
MP4 BB AB TG VNW p m=1 L=350n W=1800n
MN4 BB A  TG VPW n m=1 L=350n W=1200n

* OINV
MP5 VDD TG Y VNW p m=1 L=350n W=1800n
MN5 VSS TG Y VPW n m=1 L=350n W=1200n
.ends
