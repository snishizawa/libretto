.subckt INV_1X A YB VDD VSS VNW VPW
MP1 VDD A YB VNW p m=1 L=350n W=1800n
MN1 VSS A YB VPW n m=1 L=350n W=1200n
.ends
