.subckt AND2_1X A B Y VDD VSS VNW VPW
MP1 VDD A YB VNW p m=1    L=350n W=1800n
MP2 VDD B YB VNW p m=1    L=350n W=1800n
MN1 VSS A W1 VPW n m=1    L=350n W=1200n
MN2 W1  B YB VPW n m=1    L=350n W=1200n
MP3 VDD YB Y VNW p m=1 L=350n W=1800n
MN3 VSS YB Y VPW n m=1 L=350n W=1200n
.ends
