.subckt AOI21_1X A1 A2 B YB VDD VSS VNW VPW
MP1 VDD A1 w1  VNW p m=1 L=350n W=1800n
MP2 VDD A2 w1  VNW p m=1 L=350n W=1800n
MP3 w1  B  YB  VNW p m=1 L=350n W=1800n
MN1 VSS A1 w2  VPW n m=1 L=350n W=1200n
MN2 w2  A2 YB  VPW n m=1 L=350n W=1200n
MN3 VSS B  YB  VPW n m=1 L=350n W=1200n
.ends
