.subckt NAND3_1X A B C YB VDD VSS VNW VPW
MP1 VDD A YB  VNW p m=1 L=350n W=1800n
MP2 VDD B YB  VNW p m=1 L=350n W=1800n
MP3 VDD C YB  VNW p m=1 L=350n W=1800n
MN1 VSS A W1  VPW n m=1 L=350n W=1200n
MN2 W1  B W2  VPW n m=1 L=350n W=1200n
MN3 W2  C YB  VPW n m=1 L=350n W=1200n
.ends
