* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
X0 a_560_47# a_193_47# a_644_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_644_413# a_711_307# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_711_307# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Q a_711_307# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_465_369# a_27_47# a_560_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR a_299_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_940_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND a_711_307# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_299_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 VPWR a_711_307# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_560_47# a_27_47# a_657_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X11 VGND a_299_47# a_465_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR a_560_47# a_711_307# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_27_47# GATE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_27_47# GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 a_657_47# a_711_307# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_299_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_465_47# a_193_47# a_560_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X20 a_711_307# a_560_47# a_940_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Q a_711_307# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends
