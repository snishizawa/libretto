.subckt OA22_1X A1 A2 B Y VDD VSS VNW VPW
MP1 VDD A1 w1  VNW p m=1 L=350n W=1800n
MP2 w1  A2 YB  VNW p m=1 L=350n W=1800n
MP3 VDD B1 w2  VNW p m=1 L=350n W=1800n
MP4 w2  B2 YB  VNW p m=1 L=350n W=1800n
MN1 w3  B1 YB  VPW n m=1 L=350n W=1200n
MN2 w3  B2 YB  VPW n m=1 L=350n W=1200n
MN3 w3  A1 VSS VPW n m=1 L=350n W=1200n
MN4 w3  A2 VSS VPW n m=1 L=350n W=1200n
MP5 VDD YB Y VNW p m=1 L=350n W=1800n
MN5 VSS YB Y VPW n m=1 L=350n W=1200n
.ends
