* Library name: sg13g2_stdcell
* Cell name: sg13g2_inv_16
* View name: schematic
* Inherited view list: spectre cmos_sch cmos.sch schematic veriloga ahdl
* pspice dspf
.subckt sg13g2_inv_16 A VDD VSS Y
XX1 Y A VSS VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=16
XX0 Y A VDD VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=16
.ends
* End of subcircuit definition.
