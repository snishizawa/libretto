.subckt SEL2_1X IN0 IN1 SEL Y VDD VSS VNW VPW
* SELINV
MP1 VDD SEL SELB VNW p m=1 L=350n W=1800n
MN1 VSS SEL SELB VPW n m=1 L=350n W=1200n

* IN0INV
MP2 VDD IN0 IN0B VNW p m=1 L=350n W=1800n
MN2 VSS IN0 IN0B VPW n m=1 L=350n W=1200n

* IN1INV
MP3 VDD IN1 IN1B VNW p m=1 L=350n W=1800n
MN3 VSS IN1 IN1B VPW n m=1 L=350n W=1200n

* IN1TG
MP4 Z SELB IN1B VNW p m=1 L=350n W=1800n
MN4 Z SEL  IN1B VPW n m=1 L=350n W=1200n

* IN0TG
MP5 Z SEL  IN0B VNW p m=1 L=350n W=1800n
MN5 Z SELB IN0B VPW n m=1 L=350n W=1200n

* OUTINV
MP6 Y Z VDD VNW p m=1 L=350n W=1800n
MN6 Y Z VSS VPW n m=1 L=350n W=1200n


.ends
