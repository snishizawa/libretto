.subckt %CIRNAME% A Y VDD VSS VNW VPW
MP1 VDD A YB VNW %P% m=%MP% L=%LP%n W=%WP%n
MN1 VSS A YB VPW %N% m=%MN% L=%LN%n W=%WN%n
MP2 VDD YB Y VNW %P% m=%MP% L=%LP%n W='4*%WP%n'
MN2 VSS YB Y VPW %N% m=%MN% L=%LN%n W='4*%WN%n'
.ends
