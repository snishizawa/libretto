* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 a_86_235# A1 a_715_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND a_86_235# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_715_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND D1 a_86_235# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_86_235# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR a_86_235# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND B1 a_86_235# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR A2 a_607_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 X a_86_235# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_607_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_499_297# B1 a_607_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_86_235# D1 a_427_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_427_297# C1 a_499_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 X a_86_235# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
