* Library name: sg13g2_stdcell
* Cell name: sg13g2_sdfbbp_1
* View name: schematic
* Inherited view list: spectre cmos_sch cmos.sch schematic veriloga ahdl
* pspice dspf
.subckt sg13g2_sdfbbp_1 CLK D Q Q_N RESET_B SCD SCE SET_B VDD VSS
XX46 a_1625_93_ RESET_B VDD VDD sg13_lv_pmos w=640.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX45 a_2037_442_ a_1878_420_ a_2384_392_ VDD sg13_lv_pmos w=1.000u l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX44 VDD SET_B a_2037_442_ VDD sg13_lv_pmos w=1.000u l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX41 VDD a_622_98_ a_877_98_ VDD sg13_lv_pmos w=1.12e-06 l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX39 VDD SCE a_341_93_ VDD sg13_lv_pmos w=640.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX38 a_218_464_ D a_197_119_ VDD sg13_lv_pmos w=640.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX33 a_1092_96_ a_622_98_ a_1221_419_ VDD sg13_lv_pmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX28 a_1221_419_ a_1250_231_ VDD VDD sg13_lv_pmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX27 VDD SCE a_218_464_ VDD sg13_lv_pmos w=640.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX26 VDD a_2037_442_ Q_N VDD sg13_lv_pmos w=1.12e-06 l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX24 VDD a_1250_231_ a_1766_379_ VDD sg13_lv_pmos w=840.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX19 a_2384_392_ a_1625_93_ VDD VDD sg13_lv_pmos w=1.000u l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX17 VDD SET_B a_1250_231_ VDD sg13_lv_pmos w=840.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX16 a_27_464_ SCD VDD VDD sg13_lv_pmos w=640.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX15 a_622_98_ CLK VDD VDD sg13_lv_pmos w=1.12e-06 l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX14 a_1250_231_ a_1092_96_ a_1580_379_ VDD sg13_lv_pmos w=840.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX11 a_197_119_ a_877_98_ a_1092_96_ VDD sg13_lv_pmos w=640.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX9 a_197_119_ a_341_93_ a_27_464_ VDD sg13_lv_pmos w=640.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX8 a_2881_74_ a_2037_442_ VDD VDD sg13_lv_pmos w=840.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX7 a_1580_379_ a_1625_93_ VDD VDD sg13_lv_pmos w=840.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX6 a_1986_504_ a_2037_442_ VDD VDD sg13_lv_pmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX5 a_1878_420_ a_877_98_ a_1986_504_ VDD sg13_lv_pmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX4 a_1766_379_ a_622_98_ a_1878_420_ VDD sg13_lv_pmos w=840.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX3 VDD a_2881_74_ Q VDD sg13_lv_pmos w=1.12e-06 l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX47 a_2271_74_ a_1878_420_ a_2037_442_ VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX43 a_197_119_ a_622_98_ a_1092_96_ VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX42 a_299_119_ a_341_93_ VSS VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX40 VSS a_622_98_ a_877_98_ VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX37 a_1625_93_ RESET_B VSS VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX36 a_2061_74_ a_2037_442_ VSS VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX35 a_1418_125_ a_1092_96_ a_1250_231_ VSS sg13_lv_nmos w=550.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX34 VSS SCE a_341_93_ VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX32 VSS SET_B a_1418_125_ VSS sg13_lv_nmos w=550.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX31 a_1192_96_ a_1250_231_ VSS VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX30 a_119_119_ SCE a_197_119_ VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX29 VSS SET_B a_2271_74_ VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX25 a_1092_96_ a_877_98_ a_1192_96_ VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX23 a_197_119_ D a_299_119_ VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX22 a_2881_74_ a_2037_442_ VSS VSS sg13_lv_nmos w=550.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX21 a_1878_420_ a_622_98_ a_2061_74_ VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX20 VSS a_2881_74_ Q VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX18 VSS a_1250_231_ a_1880_119_ VSS sg13_lv_nmos w=550.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX13 a_622_98_ CLK VSS VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX12 VSS SCD a_119_119_ VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX10 a_1880_119_ a_877_98_ a_1878_420_ VSS sg13_lv_nmos w=550.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX2 a_1250_231_ a_1625_93_ a_1418_125_ VSS sg13_lv_nmos w=550.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX1 VSS a_2037_442_ Q_N VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
XX0 a_2037_442_ a_1625_93_ a_2271_74_ VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
.ends
* End of subcircuit definition.
