.subckt DFFARAS_1X CLK DATA NRST NSET Q VDD VSS VNW VPW  
*.PININFO CLK:I DATA:I NRST:I NSET:I Q:O VNW:B VPW:B
* CKB
MP11 ckb CLK VDD VNW p L=350n W=1350n
MN11 ckb CLK VSS VPW n L=350n W=900n
* CK
MP3 ck ckb VDD VNW p L=350n W=1350n
MN3 ck ckb VSS VPW n L=350n W=900n
* INCINV(D)
MP12 23 DATA VDD VNW p L=350n W=1800n
MP6 mh ck 23 VNW     p L=350n W=1800n
MN2 mh ckb 22 VPW    n L=350n W=1200n
MN12 22 DATA VSS VPW n L=350n W=1200n
* MLNAND_SETN(D)
MP15 ml NSET VDD VNW p L=350n W=1350n
MP4 ml mh VDD VNW    p L=350n W=1350n
MN4 ml mh 5 VPW      n L=350n W=900n
MN15 5 NSET VSS VPW  n L=350n W=900n
* MLNAND_RSTN(latch)
MP14 21 NRST VDD VNW p L=350n W=900n
MP7 21 ml VDD VNW    p L=350n W=900n
MN7 21 ml 8 VPW      n L=350n W=600n
MN14 8 NRST VSS VPW  n L=350n W=600n
* MLTG(latch)
MP2 mh ckb 21 VNW    p L=350n W=900n
MN6 mh ck 21 VPW     n L=350n W=600n
*TG(D)
MP1 sh ckb ml VNW p L=350n W=1350n
MN5 sh ck ml VPW  n L=350n W=900n
* SLNAND_NRST(D)
MP10 sl sh VDD VNW   p L=350n W=1350n
MP13 sl NRST VDD VNW p L=350n W=1350n
MN10 sl sh 7 VPW     n L=350n W=900n
MN13 7 NRST VSS VPW  n L=350n W=900n
* SLNAND_NSET(latch)
MP8 20 sl VDD VNW    p L=350n W=900n
MP16 20 NSET VDD VNW p L=350n W=900n
MN8 20 sl 6 VPW      n L=350n W=600n
MN16 6 NSET VSS VPW  n L=350n W=600n
* SLTG(latch)
MP5 sh ck  20 VNW     p L=350n W=900n
MN1 sh ckb 20 VPW    n L=350n W=600n

* Q(D)
MP9 Q sl VDD VNW p m=1 L=350n W=1800n
MN9 Q sl VSS VPW n m=1 L=350n W=1200n

.ENDS
