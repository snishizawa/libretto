* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__maj3_1 A B C VGND VNB VPB VPWR X
X0 a_109_341# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_265_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_27_47# B a_421_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND A a_265_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_27_47# B a_421_341# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_421_341# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_421_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_27_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_27_47# C a_109_341# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 VPWR A a_265_341# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_265_341# B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
