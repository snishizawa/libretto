* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_496_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_496_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR B1 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_926_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_672_297# A3 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_102_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_102_21# A3 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_926_297# A2 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND A1 a_496_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND A3 a_496_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR A1 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_102_21# B1 a_496_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_496_47# B1 a_102_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VGND A2 a_496_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_672_297# A2 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_496_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
